
module issp (
	source,
	probe,
	source_clk);	

	output	[31:0]	source;
	input	[63:0]	probe;
	input		source_clk;
endmodule
